module xor_gate(output c, input a, b);
    // Instantiate the built-in XOR gate primitive
    // Format: xor instance_name (output, input1, input2, ...);
    xor (c, a, b); 
endmodule
